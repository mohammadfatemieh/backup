ET@TJUETSERVER.29628:1538209710